* SPICE NETLIST
***************************************

.SUBCKT XOR2_X1 VDD A Z B VSS
** N=11 EP=5 IP=0 FDC=10
M0 2 A VSS 10 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 2 10 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 2 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 9 A Z 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 9 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 8 A 2 11 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 8 11 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 3 2 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 3 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 3 B Z 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8
** N=8 EP=8 IP=10 FDC=20
X0 1 2 3 4 5 XOR2_X1 $T=0 -1860 0 0 $X=-115 $Y=-1975
X1 1 6 7 8 5 XOR2_X1 $T=0 0 0 0 $X=-115 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=16 FDC=40
X0 1 2 4 6 8 3 5 7 ICV_1 $T=0 -3720 0 0 $X=-115 $Y=-5695
X1 1 9 11 13 8 10 12 14 ICV_1 $T=0 0 0 0 $X=-115 $Y=-1975
.ENDS
***************************************
.SUBCKT 16B_XOR VSS! VDD! a<3> a<2> a<1> a<0> O<3> O<2> O<1> O<0> b<3> b<2> b<1> b<0> a<7> a<6> a<5> a<4> O<7> O<6>
+ O<5> O<4> b<7> b<6> b<5> b<4> a<11> a<10> a<9> a<8> O<11> O<10> O<9> O<8> b<11> b<10> b<9> b<8> a<15> a<14>
+ a<13> a<12> O<15> O<14> O<13> O<12> b<15> b<14> b<13> b<12>
** N=50 EP=50 IP=56 FDC=160
X0 VDD! a<3> a<2> O<3> O<2> b<3> b<2> VSS! a<1> a<0> O<1> O<0> b<1> b<0> ICV_2 $T=-28112 297 0 90 $X=-29627 $Y=182
X1 VDD! a<7> a<6> O<7> O<6> b<7> b<6> VSS! a<5> a<4> O<5> O<4> b<5> b<4> ICV_2 $T=-20672 297 0 90 $X=-22187 $Y=182
X2 VDD! a<11> a<10> O<11> O<10> b<11> b<10> VSS! a<9> a<8> O<9> O<8> b<9> b<8> ICV_2 $T=-13232 297 0 90 $X=-14747 $Y=182
X3 VDD! a<15> a<14> O<15> O<14> b<15> b<14> VSS! a<13> a<12> O<13> O<12> b<13> b<12> ICV_2 $T=-5792 297 0 90 $X=-7307 $Y=182
.ENDS
***************************************
