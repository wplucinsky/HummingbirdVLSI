* SPICE NETLIST
***************************************

.SUBCKT SDFFR_X1 QN Q RN CK D VSS VDD
** N=31 EP=7 IP=0 FDC=42
M0 VSS 9 QN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 Q 10 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 VSS 10 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=690 $Y=215 $D=1
M3 24 RN VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=880 $Y=215 $D=1
M4 25 9 24 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.255e-14 AS=2.94e-14 PD=7.3e-07 PS=7e-07 $X=1070 $Y=215 $D=1
M5 10 11 25 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=3.255e-14 PD=7.1e-07 PS=7.3e-07 $X=1275 $Y=215 $D=1
M6 26 12 10 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=1470 $Y=215 $D=1
M7 VSS 13 26 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1660 $Y=215 $D=1
M8 11 CK VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1850 $Y=215 $D=1
M9 VSS 11 12 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.655e-14 AS=2.205e-14 PD=7.3e-07 PS=6.3e-07 $X=2190 $Y=215 $D=1
M10 27 14 VSS VSS NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.655e-14 PD=4.6e-07 PS=7.3e-07 $X=2395 $Y=320 $D=1
M11 13 12 27 VSS NMOS_VTL L=5e-08 W=9e-08 AD=2.235e-14 AS=1.26e-14 PD=7.3e-07 PS=4.6e-07 $X=2585 $Y=320 $D=1
M12 28 11 13 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.99e-14 AS=2.235e-14 PD=8e-07 PS=7.3e-07 $X=2790 $Y=215 $D=1
M13 VSS 16 28 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=3.99e-14 PD=6.3e-07 PS=8e-07 $X=3030 $Y=215 $D=1
M14 29 13 14 VSS NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=9.45e-15 PD=4.6e-07 PS=3.9e-07 $X=3370 $Y=215 $D=1
M15 VSS RN 29 VSS NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.26e-14 PD=7e-07 PS=4.6e-07 $X=3560 $Y=215 $D=1
M16 30 SI VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.1e-14 PD=7e-07 PS=7e-07 $X=3750 $Y=215 $D=1
M17 16 SE 30 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.94e-14 PD=9.5e-07 PS=7e-07 $X=3940 $Y=215 $D=1
M18 31 18 16 VSS NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=9.5e-07 $X=4130 $Y=90 $D=1
M19 VSS D 31 VSS NMOS_VTL L=5e-08 W=2.75e-07 AD=3.395e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=4320 $Y=90 $D=1
M20 18 SE VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=3.395e-14 PD=6.3e-07 PS=8.3e-07 $X=4510 $Y=155 $D=1
M21 VDD 9 QN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M22 Q 10 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M23 VDD 10 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=690 $Y=995 $D=0
M24 8 RN VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=880 $Y=995 $D=0
M25 VDD 9 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1070 $Y=995 $D=0
M26 10 12 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1410 $Y=815 $D=0
M27 19 11 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1600 $Y=815 $D=0
M28 VDD 13 19 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1790 $Y=815 $D=0
M29 11 CK VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1980 $Y=815 $D=0
M30 VDD 11 12 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=2320 $Y=870 $D=0
M31 20 14 VDD VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=2510 $Y=1010 $D=0
M32 13 11 20 VDD PMOS_VTL L=5e-08 W=9e-08 AD=4.815e-14 AS=1.26e-14 PD=1.1e-06 PS=4.6e-07 $X=2700 $Y=1010 $D=0
M33 21 12 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.815e-14 PD=9.1e-07 PS=1.1e-06 $X=2985 $Y=870 $D=0
M34 VDD 16 21 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.88e-14 AS=4.41e-14 PD=9.2e-07 PS=9.1e-07 $X=3175 $Y=870 $D=0
M35 14 13 VDD VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.88e-14 PD=4.6e-07 PS=9.2e-07 $X=3370 $Y=1095 $D=0
M36 VDD RN 14 VDD PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.26e-14 PD=9.1e-07 PS=4.6e-07 $X=3560 $Y=1095 $D=0
M37 22 SI VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=2.835e-14 PD=9.1e-07 PS=9.1e-07 $X=3750 $Y=870 $D=0
M38 16 18 22 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=4.41e-14 PD=1.12e-06 PS=9.1e-07 $X=3940 $Y=870 $D=0
M39 23 SE 16 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=4130 $Y=870 $D=0
M40 VDD D 23 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.145e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=4320 $Y=870 $D=0
M41 18 SE VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=5.145e-14 PD=8.4e-07 PS=1.12e-06 $X=4510 $Y=975 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=14 FDC=84
X0 3 4 5 6 7 1 2 SDFFR_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 8 9 5 6 10 1 2 SDFFR_X1 $T=4746 0 0 0 $X=4631 $Y=-115
.ENDS
***************************************
.SUBCKT 16_bit_register RN CK QN<0> VDD! VSS! Q<0> D<0> QN<1> Q<1> D<1> QN<2> Q<2> D<2> QN<3> Q<3> D<3> QN<4> Q<4> D<4> QN<5>
+ Q<5> D<5> QN<6> Q<6> D<6> QN<7> Q<7> D<7> QN<8> Q<8> D<8> QN<9> Q<9> D<9> QN<10> Q<10> D<10> QN<11> Q<11> D<11>
+ QN<12> Q<12> D<12> QN<13> Q<13> D<13> QN<14> Q<14> D<14> QN<15> Q<15> D<15>
** N=52 EP=52 IP=92 FDC=672
X0 QN<8> Q<8> RN CK D<8> VSS! VDD! SDFFR_X1 $T=41619 441 0 0 $X=41504 $Y=326
X1 QN<9> Q<9> RN CK D<9> VSS! VDD! SDFFR_X1 $T=46368 441 0 0 $X=46253 $Y=326
X2 QN<12> Q<12> RN CK D<12> VSS! VDD! SDFFR_X1 $T=60600 441 0 0 $X=60485 $Y=326
X3 QN<13> Q<13> RN CK D<13> VSS! VDD! SDFFR_X1 $T=65343 441 0 0 $X=65228 $Y=326
X4 QN<14> Q<14> RN CK D<14> VSS! VDD! SDFFR_X1 $T=70092 441 0 0 $X=69977 $Y=326
X5 QN<15> Q<15> RN CK D<15> VSS! VDD! SDFFR_X1 $T=74829 441 0 0 $X=74714 $Y=326
X6 VSS! VDD! QN<0> Q<0> RN CK D<0> QN<1> Q<1> D<1> ICV_1 $T=3657 441 0 0 $X=3542 $Y=326
X7 VSS! VDD! QN<2> Q<2> RN CK D<2> QN<3> Q<3> D<3> ICV_1 $T=13149 441 0 0 $X=13034 $Y=326
X8 VSS! VDD! QN<4> Q<4> RN CK D<4> QN<5> Q<5> D<5> ICV_1 $T=22635 441 0 0 $X=22520 $Y=326
X9 VSS! VDD! QN<6> Q<6> RN CK D<6> QN<7> Q<7> D<7> ICV_1 $T=32127 441 0 0 $X=32012 $Y=326
X10 VSS! VDD! QN<10> Q<10> RN CK D<10> QN<11> Q<11> D<11> ICV_1 $T=51108 441 0 0 $X=50993 $Y=326
.ENDS
***************************************
