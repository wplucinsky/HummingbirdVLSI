* SPICE NETLIST
***************************************

.SUBCKT AND2_X1 A1 A2 VSS VDD ZN
** N=9 EP=5 IP=0 FDC=6
M0 7 A1 6 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 7 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 6 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 6 A1 VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 6 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 6 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS
** N=11 EP=5 IP=0 FDC=10
M0 6 A VSS 10 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 6 10 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 6 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 9 A Z 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 9 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 8 A 6 11 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 8 11 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 7 6 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 7 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 7 B Z 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FullAdder A B Cin Cout VSS! VDD! Sum
** N=14 EP=7 IP=20 FDC=38
M0 11 8 VSS! 13 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=337 $Y=-1566 $D=1
M1 VSS! 9 11 13 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=527 $Y=-1566 $D=1
M2 Cout 11 VSS! 13 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=717 $Y=-1566 $D=1
M3 12 8 11 14 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=337 $Y=-661 $D=0
M4 VDD! 9 12 14 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=527 $Y=-661 $D=0
M5 Cout 11 VDD! 14 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=717 $Y=-976 $D=0
X6 A B VSS! VDD! 9 AND2_X1 $T=2547 -1683 0 0 $X=2432 $Y=-1798
X7 Cin 10 VSS! VDD! 8 AND2_X1 $T=6975 -1683 0 0 $X=6860 $Y=-1798
X8 VDD! A 10 B VSS! XOR2_X1 $T=4788 -1683 0 0 $X=4673 $Y=-1798
X9 VDD! 10 Sum Cin VSS! XOR2_X1 $T=9663 -1683 0 0 $X=9548 $Y=-1798
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8 9 10 11
** N=13 EP=11 IP=14 FDC=76
X0 7 8 3 1 12 13 2 FullAdder $T=0 0 0 0 $X=77 $Y=-2229
X1 9 10 11 3 4 5 6 FullAdder $T=11892 0 0 0 $X=11969 $Y=-2229
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19
** N=21 EP=19 IP=22 FDC=152
X0 1 2 3 20 21 4 11 12 13 14 5 ICV_1 $T=0 0 0 0 $X=77 $Y=-2229
X1 5 6 7 8 9 10 15 16 17 18 19 ICV_1 $T=23790 0 0 0 $X=23867 $Y=-2229
.ENDS
***************************************
.SUBCKT 16BitAdder cout VSS! VDD! sum<15> sum<14> sum<13> sum<12> sum<11> sum<10> sum<9> sum<8> sum<7> sum<6> sum<5> sum<4> sum<3> sum<2> sum<1> sum<0> A<15>
+ B<15> A<14> B<14> A<13> B<13> A<12> B<12> A<11> B<11> A<10> B<10> A<9> B<9> A<8> B<8> A<7> B<7> A<6> B<6> A<5>
+ B<5> A<4> B<4> A<3> B<3> A<2> B<2> A<1> B<1> A<0> B<0> GND!
** N=73 EP=52 IP=76 FDC=608
X0 cout sum<15> 2 sum<14> 3 sum<13> 4 22 23 sum<12> A<15> B<15> A<14> B<14> A<13> B<13> A<12> B<12> 5 ICV_2 $T=2265 -1812 0 0 $X=2342 $Y=-4041
X1 5 sum<11> 6 sum<10> 7 sum<9> 8 28 29 sum<8> A<11> B<11> A<10> B<10> A<9> B<9> A<8> B<8> 9 ICV_2 $T=49956 -1812 0 0 $X=50033 $Y=-4041
X2 9 sum<7> 10 sum<6> 11 sum<5> 12 34 35 sum<4> A<7> B<7> A<6> B<6> A<5> B<5> A<4> B<4> 13 ICV_2 $T=97527 -1812 0 0 $X=97604 $Y=-4041
X3 13 sum<3> 14 sum<2> 15 sum<1> 16 VSS! VDD! sum<0> A<3> B<3> A<2> B<2> A<1> B<1> A<0> B<0> GND! ICV_2 $T=145110 -1812 0 0 $X=145187 $Y=-4041
.ENDS
***************************************
