* SPICE NETLIST
***************************************

.SUBCKT dff 1 2 3 4 5 a b 8 9 10 Out 12 13 14 gnd! 16 17 vdd!
** N=28 EP=18 IP=0 FDC=32
M0 21 a gnd! gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.8e-14 AS=2.1e-14 PD=6.8e-07 PS=6.1e-07 $X=-3830 $Y=405 $D=3
M1 1 2 21 gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.2e-14 AS=2.8e-14 PD=6.2e-07 PS=6.8e-07 $X=-3450 $Y=405 $D=3
M2 22 1 gnd! gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.8e-14 AS=2.1e-14 PD=6.8e-07 PS=6.1e-07 $X=-2325 $Y=300 $D=3
M3 2 b 22 gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.2e-14 AS=2.8e-14 PD=6.2e-07 PS=6.8e-07 $X=-1945 $Y=300 $D=3
M4 23 2 gnd! gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.8e-14 AS=2.1e-14 PD=6.8e-07 PS=6.1e-07 $X=-825 $Y=405 $D=3
M5 9 8 23 gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.2e-14 AS=2.8e-14 PD=6.2e-07 PS=6.8e-07 $X=-445 $Y=405 $D=3
M6 24 9 gnd! gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.8e-14 AS=2.1e-14 PD=6.8e-07 PS=6.1e-07 $X=685 $Y=405 $D=3
M7 10 3 24 gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.2e-14 AS=2.8e-14 PD=6.2e-07 PS=6.8e-07 $X=1065 $Y=405 $D=3
M8 25 10 gnd! gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.8e-14 AS=2.1e-14 PD=6.8e-07 PS=6.1e-07 $X=2180 $Y=405 $D=3
M9 Out 13 25 gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.2e-14 AS=2.8e-14 PD=6.2e-07 PS=6.8e-07 $X=2560 $Y=405 $D=3
M10 26 12 gnd! gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.8e-14 AS=2.1e-14 PD=6.8e-07 PS=6.1e-07 $X=3685 $Y=405 $D=3
M11 13 4 26 gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.2e-14 AS=2.8e-14 PD=6.2e-07 PS=6.8e-07 $X=4065 $Y=405 $D=3
M12 27 4 gnd! gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.8e-14 AS=2.1e-14 PD=6.8e-07 PS=6.1e-07 $X=5170 $Y=405 $D=3
M13 14 17 27 gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.2e-14 AS=2.8e-14 PD=6.2e-07 PS=6.8e-07 $X=5550 $Y=405 $D=3
M14 28 5 gnd! gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.8e-14 AS=2.1e-14 PD=6.8e-07 PS=6.1e-07 $X=6675 $Y=405 $D=3
M15 17 16 28 gnd! NMOS_VTH L=5e-08 W=2e-07 AD=2.2e-14 AS=2.8e-14 PD=6.2e-07 PS=6.8e-07 $X=7055 $Y=405 $D=3
M16 1 a vdd! vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.835e-14 AS=2.12625e-14 PD=6.85e-07 PS=6.15e-07 $X=-3830 $Y=1770 $D=2
M17 vdd! 2 1 vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.2275e-14 AS=2.835e-14 PD=6.25e-07 PS=6.85e-07 $X=-3450 $Y=1770 $D=2
M18 2 1 vdd! vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.835e-14 AS=2.12625e-14 PD=6.85e-07 PS=6.15e-07 $X=-2325 $Y=1770 $D=2
M19 vdd! b 2 vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.2275e-14 AS=2.835e-14 PD=6.25e-07 PS=6.85e-07 $X=-1945 $Y=1770 $D=2
M20 9 2 vdd! vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.835e-14 AS=2.12625e-14 PD=6.85e-07 PS=6.15e-07 $X=-825 $Y=1770 $D=2
M21 vdd! 8 9 vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.2275e-14 AS=2.835e-14 PD=6.25e-07 PS=6.85e-07 $X=-445 $Y=1770 $D=2
M22 10 9 vdd! vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.835e-14 AS=2.12625e-14 PD=6.85e-07 PS=6.15e-07 $X=685 $Y=1770 $D=2
M23 vdd! 3 10 vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.2275e-14 AS=2.835e-14 PD=6.25e-07 PS=6.85e-07 $X=1065 $Y=1770 $D=2
M24 Out 10 vdd! vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.835e-14 AS=2.12625e-14 PD=6.85e-07 PS=6.15e-07 $X=2180 $Y=1770 $D=2
M25 vdd! 13 Out vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.2275e-14 AS=2.835e-14 PD=6.25e-07 PS=6.85e-07 $X=2560 $Y=1770 $D=2
M26 13 12 vdd! vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.835e-14 AS=2.12625e-14 PD=6.85e-07 PS=6.15e-07 $X=3685 $Y=1770 $D=2
M27 vdd! 4 13 vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.2275e-14 AS=2.835e-14 PD=6.25e-07 PS=6.85e-07 $X=4065 $Y=1770 $D=2
M28 14 4 vdd! vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.835e-14 AS=2.12625e-14 PD=6.85e-07 PS=6.15e-07 $X=5170 $Y=1770 $D=2
M29 vdd! 17 14 vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.2275e-14 AS=2.835e-14 PD=6.25e-07 PS=6.85e-07 $X=5550 $Y=1770 $D=2
M30 17 5 vdd! vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.835e-14 AS=2.12625e-14 PD=6.85e-07 PS=6.15e-07 $X=6675 $Y=1770 $D=2
M31 vdd! 16 17 vdd! PMOS_VTH L=5e-08 W=2.025e-07 AD=2.2275e-14 AS=2.835e-14 PD=6.25e-07 PS=6.85e-07 $X=7055 $Y=1770 $D=2
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
