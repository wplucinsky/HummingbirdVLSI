* SPICE NETLIST
***************************************

.SUBCKT DFFR_X1 D VSS VDD Q
** N=25 EP=4 IP=0 FDC=32
M0 VSS CK 5 24 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=140 $D=1
M1 10 5 VSS 24 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=335 $Y=140 $D=1
M2 18 D VSS 24 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=2.8875e-14 PD=8.3e-07 PS=7.6e-07 $X=675 $Y=215 $D=1
M3 7 5 18 24 NMOS_VTL L=5e-08 W=2.75e-07 AD=2.555e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=865 $Y=215 $D=1
M4 19 10 7 24 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.555e-14 PD=4.6e-07 PS=8.3e-07 $X=1055 $Y=305 $D=1
M5 20 9 19 24 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1245 $Y=305 $D=1
M6 VSS RN 20 24 NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14 PD=3.9e-07 PS=4.6e-07 $X=1435 $Y=305 $D=1
M7 VSS 7 9 24 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.41e-14 AS=2.205e-14 PD=8.4e-07 PS=6.3e-07 $X=1790 $Y=215 $D=1
M8 21 7 VSS 24 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.41e-14 PD=7e-07 PS=8.4e-07 $X=2050 $Y=215 $D=1
M9 12 10 21 24 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2240 $Y=215 $D=1
M10 22 5 12 24 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=2430 $Y=215 $D=1
M11 VSS 14 22 24 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.26e-14 PD=7e-07 PS=4.6e-07 $X=2620 $Y=215 $D=1
M12 23 RN VSS 24 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.1e-14 PD=7e-07 PS=7e-07 $X=2810 $Y=215 $D=1
M13 14 12 23 24 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=3000 $Y=215 $D=1
M14 VSS 12 QN 24 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=3385 $Y=90 $D=1
M15 Q 14 VSS 24 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=3575 $Y=90 $D=1
M16 VDD CK 5 25 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M17 10 5 VDD 25 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M18 15 D VDD 25 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=4.41e-14 PD=1.12e-06 PS=1.05e-06 $X=675 $Y=840 $D=0
M19 7 10 15 25 PMOS_VTL L=5e-08 W=4.2e-07 AD=3.57e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=865 $Y=840 $D=0
M20 8 5 7 25 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.57e-14 PD=4.6e-07 PS=1.12e-06 $X=1055 $Y=1020 $D=0
M21 VDD 9 8 25 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1245 $Y=1020 $D=0
M22 8 RN VDD 25 PMOS_VTL L=5e-08 W=9e-08 AD=1.035e-14 AS=1.26e-14 PD=4.1e-07 PS=4.6e-07 $X=1435 $Y=1020 $D=0
M23 VDD 7 9 25 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.465e-14 PD=1.05e-06 PS=8.5e-07 $X=1790 $Y=855 $D=0
M24 16 7 VDD 25 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.05e-06 $X=2050 $Y=855 $D=0
M25 12 5 16 25 PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2240 $Y=855 $D=0
M26 17 10 12 25 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=2430 $Y=995 $D=0
M27 VDD 14 17 25 PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.26e-14 PD=9.1e-07 PS=4.6e-07 $X=2620 $Y=995 $D=0
M28 14 RN VDD 25 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=2.835e-14 PD=9.1e-07 PS=9.1e-07 $X=2810 $Y=995 $D=0
M29 VDD 12 14 25 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=3000 $Y=995 $D=0
M30 VDD 12 QN 25 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=3385 $Y=680 $D=0
M31 Q 14 VDD 25 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3575 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5
** N=5 EP=5 IP=8 FDC=64
X0 3 1 2 4 DFFR_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 4 1 2 5 DFFR_X1 $T=4255 0 0 0 $X=4140 $Y=-115
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7
** N=7 EP=7 IP=10 FDC=128
X0 1 2 3 4 5 ICV_1 $T=0 0 0 0 $X=-115 $Y=-115
X1 1 2 5 6 7 ICV_1 $T=8510 0 0 0 $X=8395 $Y=-115
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS
** N=11 EP=5 IP=0 FDC=10
M0 6 A VSS 10 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 6 10 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 6 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 9 A Z 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 9 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 8 A 6 11 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 8 11 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 7 6 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 7 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 7 B Z 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT LFSR Out<15> Out<0> Out<14> Out<13> Out<12> Out<11> Out<10> Out<9> Out<8> Out<7> Out<6> Out<5> Out<4> Out<3> Out<2> Out<1> VSS! VDD!
** N=22 EP=18 IP=55 FDC=542
X0 22 VSS! VDD! Out<15> DFFR_X1 $T=-105 185 0 0 $X=-220 $Y=70
X1 Out<15> VSS! VDD! 2 DFFR_X1 $T=4210 185 0 0 $X=4095 $Y=70
X2 Out<14> VSS! VDD! 5 DFFR_X1 $T=10060 185 0 0 $X=9945 $Y=70
X3 Out<1> VSS! VDD! Out<0> DFFR_X1 $T=68570 185 0 0 $X=68455 $Y=70
X4 VSS! VDD! Out<13> Out<12> 8 ICV_1 $T=15910 185 0 0 $X=15795 $Y=70
X5 VSS! VDD! Out<3> Out<2> Out<1> ICV_1 $T=60055 185 0 0 $X=59940 $Y=70
X6 VSS! VDD! Out<11> Out<10> Out<9> Out<8> Out<7> ICV_2 $T=26015 185 0 0 $X=25900 $Y=70
X7 VSS! VDD! Out<7> Out<6> Out<5> Out<4> Out<3> ICV_2 $T=43035 185 0 0 $X=42920 $Y=70
X8 VDD! 2 Out<14> Out<0> VSS! XOR2_X1 $T=8465 185 0 0 $X=8350 $Y=70
X9 VDD! 5 Out<13> Out<0> VSS! XOR2_X1 $T=14315 185 0 0 $X=14200 $Y=70
X10 VDD! 8 Out<11> Out<0> VSS! XOR2_X1 $T=24420 185 0 0 $X=24305 $Y=70
.ENDS
***************************************
