* SPICE NETLIST
***************************************

.SUBCKT INV_X1 A VSS VDD ZN 5 6
** N=6 EP=6 IP=0 FDC=2
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN
** N=9 EP=5 IP=0 FDC=6
M0 7 A1 3 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 7 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 3 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 3 A1 VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 3 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 3 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT 2x4_decoder A0 A1 VSS! VDD! D<0> D<1> D<2> D<3>
** N=12 EP=8 IP=32 FDC=28
X0 A0 VSS! VDD! 2 VSS! VDD! INV_X1 $T=1482 462 0 0 $X=1367 $Y=347
X1 A1 VSS! VDD! 4 11 12 INV_X1 $T=2433 462 0 0 $X=2318 $Y=347
X2 4 2 VSS! VDD! D<0> AND2_X1 $T=3579 462 0 0 $X=3464 $Y=347
X3 A0 4 VSS! VDD! D<1> AND2_X1 $T=5247 462 0 0 $X=5132 $Y=347
X4 A1 2 VSS! VDD! D<2> AND2_X1 $T=6906 462 0 0 $X=6791 $Y=347
X5 A0 A1 VSS! VDD! D<3> AND2_X1 $T=8469 462 0 0 $X=8354 $Y=347
.ENDS
***************************************
