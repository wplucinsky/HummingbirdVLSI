* SPICE NETLIST
***************************************

.SUBCKT XOR2_X1 VDD A Z B VSS
** N=11 EP=5 IP=0 FDC=10
M0 2 A VSS 10 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 2 10 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 2 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 9 A Z 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 9 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 8 A 2 11 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 8 11 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 3 2 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 3 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 3 B Z 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT 3i_XOR VSS! VDD! A B out C
** N=7 EP=6 IP=10 FDC=20
X0 VDD! A 1 B VSS! XOR2_X1 $T=-5760 801 0 0 $X=-5875 $Y=686
X1 VDD! 1 out C VSS! XOR2_X1 $T=-3471 801 0 0 $X=-3586 $Y=686
.ENDS
***************************************
.SUBCKT ICV_1 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 IP=12 FDC=40
X0 1 2 3 4 6 5 3i_XOR $T=0 0 0 0 $X=-5875 $Y=686
X1 1 2 7 8 10 9 3i_XOR $T=4677 0 0 0 $X=-1198 $Y=686
.ENDS
***************************************
.SUBCKT ICV_2 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18
** N=18 EP=18 IP=20 FDC=80
X0 1 2 3 4 5 6 7 8 9 10 ICV_1 $T=0 0 0 0 $X=-5875 $Y=686
X1 1 2 11 12 13 14 15 16 17 18 ICV_1 $T=9327 0 0 0 $X=3452 $Y=686
.ENDS
***************************************
.SUBCKT LTB m<5> m<8> m<4> m<7> m<3> m<6> m<2> m<1> GND! m<15> O<15> m<14> O<14> m<13> O<13> m<12> O<12> m<11> O<11> m<10>
+ O<10> O<9> O<8> O<7> O<6> O<5> O<4> O<3> O<2> O<1> O<0>
** N=35 EP=31 IP=72 FDC=320
X0 12 13 m<15> 1 m<5> O<15> m<14> m<8> m<4> O<14> m<13> m<7> m<3> O<13> m<12> m<6> m<2> O<12> ICV_2 $T=6951 -3267 0 0 $X=1076 $Y=-2581
X1 12 13 m<11> m<5> m<1> O<11> m<10> m<4> 10 O<10> 1 m<3> GND! O<9> m<8> m<2> GND! O<8> ICV_2 $T=25527 -3267 0 0 $X=19652 $Y=-2581
X2 12 13 m<7> m<1> GND! O<7> m<6> 10 GND! O<6> m<5> GND! GND! O<5> m<4> GND! GND! O<4> ICV_2 $T=44088 -3267 0 0 $X=38213 $Y=-2581
X3 12 13 m<3> GND! GND! O<3> m<2> GND! GND! O<2> m<1> GND! GND! O<1> 10 GND! GND! O<0> ICV_2 $T=62664 -3267 0 0 $X=56789 $Y=-2581
.ENDS
***************************************
